library verilog;
use verilog.vl_types.all;
entity FloatingPointAdder_vlg_vec_tst is
end FloatingPointAdder_vlg_vec_tst;
