library ieee;
use ieee.std_logic_1164.all;

entity HalfAdder is
	port(
		a, b : in std_logic;
		s, c : out std_logic
	);
	end HalfAdder;

architecture rtl of HalfAdder is 
	begin
		c <= a and b;
		s <= a xor b;

end rtl;

