library verilog;
use verilog.vl_types.all;
entity AdderDataPath_vlg_vec_tst is
end AdderDataPath_vlg_vec_tst;
