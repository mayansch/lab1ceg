library verilog;
use verilog.vl_types.all;
entity FloatingPointMultiplier_vlg_vec_tst is
end FloatingPointMultiplier_vlg_vec_tst;
